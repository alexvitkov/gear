inc := x => x + 1;
add2 := x => inc(inc(x));
